LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY BCDCount2 IS
	PORT (Clear,Enable,Clock: IN STD_LOGIC;
			BCD_0, BCD_1: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END BCDCount2;

ARCHITECTURE BEHAVIOUR OF BCDCount2 IS

SIGNAL OR_0, OR_1, AND_0, AND_1: STD_LOGIC; --X = output from XOR gates, M = output from MUX gates
SIGNAL D, Q0, Q1: STD_LOGIC_VECTOR(3 DOWNTO 0);  -- A = output of AND gates

BEGIN
D <= "0000";
OR_0 <= Clear OR AND_0;
OR_1 <= Clear OR AND_1;
step1: ENTITY WORK.Count4 PORT MAP(OR_0,Enable,Clock,D,Q0);
AND_0 <= Q0(0) AND Q0(3);
step2: ENTITY WORK.Count4 PORT MAP(OR_1,AND_0,Clock,D,Q1);
AND_1 <= Q1(0) AND Q1(3) AND AND_0;
BCD_0 <= Q0;
BCD_1 <= Q1;
END BEHAVIOUR;